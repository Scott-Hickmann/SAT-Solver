module k(
  input wire s,
  input wire c,
  output reg 
);